module and_gate(O,A,B);
  input A,B;
  output O;
  and(O,A,B);
endmodule